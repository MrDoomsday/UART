//---------------------------------------------------------------------------------------
// uart receive module  
//
//---------------------------------------------------------------------------------------

module uart_rx 
(
// modules inputs and outputs 
	input 			clock,			// global clock input 
	input 			reset,			// global reset input 

	input 			pbit,			// enable parity bit
	input 			ptype,			// type parity bit, 0 - even, 1 - odd
	input 	[1:0] 	sbit,			// count stop bit, 2'b00 - 1 stop bit, 2'b01 - 2 stop bit, 2'b10 - 3 stop bit, 2'b11 - 3 stop bit;
	
	input				ce_8,			// baud rate multiplyed by 16 - generated by baud module 
	input				ser_in,			// serial data input 
	output	reg [7:0]	rx_data,		// data byte received 
	output 	reg			new_rx_data,	// signs that a new byte was received 
	output 	reg			pbit_error
);
//---------------------------------------------------------------------------------------


// internal wires 
wire ce_1;		// clock enable at bit rate 
wire ce_1_mid;	// clock enable at the middle of each bit - used to sample data 

// internal registers 
reg [1:0] in_sync;
reg rx_busy; 
reg [2:0]	count8;
reg [3:0]	bit_count;
reg [8:0]	data_buf;
reg 		pbit_r;
reg 		ptype_r;
reg [1:0] 	sbit_r;
//---------------------------------------------------------------------------------------
// module implementation 
// input async input is sampled twice 
always @ (posedge clock or posedge reset) begin 
	if (reset) in_sync <= 2'b11;
	else in_sync <= {in_sync[0], ser_in};
end 

// a counter to count 16 pulses of ce_8 to generate the ce_1 and ce_1_mid pulses.
// this counter is used to detect the start bit while the receiver is not receiving and 
// signs the sampling cycle during reception. 
always @ (posedge clock or posedge reset) begin
	if (reset) count8 <= 3'b0;
	else if (ce_8) begin 
		if (rx_busy | (in_sync[1] == 1'b0)) count8 <= count8 + 3'b1;
		else count8 <= 3'b0;
	end 
end 

// ce_1 pulse indicating expected end of current bit 
assign ce_1 = (count8 == 3'b111) & ce_8;
// ce_1_mid pulse indication the sampling clock cycle of the current data bit 
assign ce_1_mid = (count8 == 3'b011) & ce_8;

// receiving busy flag and capture control bits
always @ (posedge clock or posedge reset) begin 
	if (reset) begin 
		rx_busy <= 1'b0;
		pbit_r 	<= 1'b0;
		ptype_r <= 1'b0;
		sbit_r 	<= 2'b00;
	end
	else if (~rx_busy & ce_1_mid) begin
		rx_busy <= 1'b1;
		pbit_r <= pbit;
		ptype_r <= ptype;
		sbit_r <= sbit;
	end
	else if (rx_busy & (bit_count == (4'h8 + {2'b000, pbit_r})) & ce_1_mid) rx_busy <= 1'b0;
end 

// bit counter 
always @ (posedge clock or posedge reset) begin 
	if (reset) bit_count <= 4'h0;
	else if (~rx_busy) bit_count <= 4'h0;
	else if (rx_busy & ce_1_mid) bit_count <= bit_count + 4'h1;
end

// data buffer shift register 
always @ (posedge clock or posedge reset) begin 
	if (reset) data_buf <= 9'h0;
	else if (rx_busy & ce_1_mid) data_buf <= {in_sync[1], data_buf[8:1]};
end

// data output and flag 
wire parity_check = ^data_buf[7:0] == data_buf[8];

always @ (posedge clock or posedge reset) begin 
	if (reset) begin 
		rx_data <= 8'h0;
		new_rx_data <= 1'b0;
		pbit_error <= 1'b0;
	end 
	else if (rx_busy & (bit_count == (4'h8 + {2'b000, pbit_r})) & ce_1) begin 
		rx_data <= pbit_r ? data_buf[7:0] : data_buf[8:1];
		new_rx_data <= 1'b1;
		pbit_error <= pbit_r & (ptype_r ? parity_check : ~parity_check);
	end 
	else new_rx_data <= 1'b0;
end

endmodule
//---------------------------------------------------------------------------------------
//						Th.. Th.. Th.. Thats all folks !!!
//---------------------------------------------------------------------------------------
