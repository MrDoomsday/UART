//---------------------------------------------------------------------------------------
// uart transmit module  
//
//---------------------------------------------------------------------------------------

module uart_tx  
(
	//---------------------------------------------------------------------------------------
	// modules inputs and outputs 
	input 			clock,			// global clock input 
	input 			reset,			// global reset input 

	input 			pbit,			// enable parity bit
	input 			ptype,			// type parity bit, 0 - even, 1 - odd
	input 	[1:0] 	sbit,			// count stop bit, 2'b00 - 1 stop bit, 2'b01 - 2 stop bit, 2'b10 - 3 stop bit, 2'b11 - 3 stop bit;

	input			ce_8,			// baud rate multiplyed by 16 - generated by baud module 
	input	[7:0]	tx_data,		// data byte to transmit 
	input			new_tx_data,	// asserted to indicate that there is a new data byte for transmission 
	output	reg		ser_out,		// serial data output 
	output 	reg		tx_busy			// signs that transmitter is busy 
);


// internal wires 
wire ce_1;		// clock enable at bit rate 

// internal registers 
reg [2:0]	count8;
reg [3:0]	bit_count;
reg [9:0]	data_buf;
reg 		pbit_r;
reg 		ptype_r;
wire 		parity_bit;
reg [1:0] 	sbit_r;
//---------------------------------------------------------------------------------------
// module implementation 
// a counter to count 16 pulses of ce_8 to generate the ce_1 pulse 
always @ (posedge clock or posedge reset) begin
	if (reset)  count8 <= 3'b0;
	else if (tx_busy & ce_8) count8 <= count8 + 3'b1;
	else if (~tx_busy) count8 <= 3'b0;
end 

// ce_1 pulse indicating output data bit should be updated 
assign ce_1 = (count8 == 3'b111) & ce_8;

// tx_busy flag and capture control bits
always @ (posedge clock or posedge reset) begin
	if (reset) begin 
		tx_busy <= 1'b0;
		pbit_r 	<= 1'b0;
		ptype_r <= 1'b0;
		sbit_r 	<= 2'b00;
	end
	else if (~tx_busy & new_tx_data) begin
		tx_busy <= 1'b1;
		pbit_r <= pbit;
		ptype_r<= ptype;
		sbit_r <= sbit;
	end
	else if (tx_busy & (bit_count == 4'(4'h9 + {3'b000, pbit_r} + {2'b00, sbit_r})) & ce_1) tx_busy <= 1'b0;
end 

assign parity_bit = ^tx_data;

// output bit counter 
always @ (posedge clock or posedge reset) begin
	if (reset) bit_count <= 4'h0;
	else if (tx_busy & ce_1) bit_count <= bit_count + 4'h1;
	else if (~tx_busy) bit_count <= 4'h0;
end 

// data shift register 
always @ (posedge clock or posedge reset) begin
	if (reset) data_buf <= 9'b0;
	else if (~tx_busy) data_buf <= {(pbit ? (ptype ? ~parity_bit : parity_bit) : 1'b1), tx_data, 1'b0}; // add check bit
	else if (tx_busy & ce_1) data_buf <= {1'b1, data_buf[9:1]};
end 

// output data bit 
always @ (posedge clock or posedge reset) begin
	if (reset) ser_out <= 1'b1;
	else if (tx_busy) ser_out <= data_buf[0];
	else ser_out <= 1'b1;
end 

endmodule
//---------------------------------------------------------------------------------------
//						Th.. Th.. Th.. Thats all folks !!!
//---------------------------------------------------------------------------------------