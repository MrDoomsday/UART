module uart_rx_tx (
    input clk,
    input reset_n,

    //tx data
    input   bit     [7:0]   tx_data_i,
    input   bit             tx_valid_i,
    output  bit             tx_ready_o,

    //rx data
    output  bit     [7:0]   rx_data_o,
    output  bit             rx_pbit_error,
    output  bit             rx_valid_o,


    input   bit     uart_rx,
    output  bit     uart_tx,

    //control register
    input   bit             cr_pbit, // enable parity bit
    input   bit     [1:0]   cr_sbit, // count stop bit, 2'b00 - 1 stop bit, 2'b01 - 2 stop bit, 2'b10 - 3 stop bit, 2'b11 - 3 stop bit;
	input 	bit				cr_ptype,// type parity bit, 0 - even, 1 - odd
    input   bit     [15:0]  cr_baud_freq,
    input   bit     [15:0]	cr_baud_limit

);

/***********************************************************************************************************************/
/***********************************************************************************************************************/
/*******************************************        DECLARATION         ************************************************/
/***********************************************************************************************************************/
/***********************************************************************************************************************/
wire ce_16;
wire tx_busy;

/***********************************************************************************************************************/
/***********************************************************************************************************************/
/*******************************************           INSTANCE          ***********************************************/
/***********************************************************************************************************************/
/***********************************************************************************************************************/

baud_gen baud_gen_inst(
	//---------------------------------------------------------------------------------------
	// modules inputs and outputs 
	.clock      (clk),		// global clock input 
	.reset      (~reset_n),		// global reset input 
	.ce_16      (ce_16),		// baud rate multiplyed by 16 
	.baud_freq  (cr_baud_freq),	// baud rate setting registers - see header description 
	.baud_limit (cr_baud_limit)
);



uart_tx uart_tx_inst (
	//---------------------------------------------------------------------------------------
	// modules inputs and outputs 
	.clock      (clk),			// global clock input 
	.reset      (~reset_n),			// global reset input 

	.pbit       (cr_pbit),			// enable parity bit
	.ptype		(cr_ptype),			// type parity bit, 0 - even, 1 - odd
	.sbit       (cr_sbit),			// count stop bit, 2'b00 - 1 stop bit, 2'b01 - 2 stop bit, 2'b10 - 3 stop bit, 2'b11 - 3 stop bit;

	.ce_16      (ce_16),			// baud rate multiplyed by 16 - generated by baud module 
	.tx_data    (tx_data_i),		// data byte to transmit 
	.new_tx_data(tx_valid_i),	// asserted to indicate that there is a new data byte for transmission 
	.ser_out    (uart_tx),		// serial data output 
	.tx_busy    (tx_busy)		// signs that transmitter is busy 
);

assign tx_ready_o = ~tx_busy;


uart_rx uart_rx_inst(
// modules inputs and outputs 
	.clock      (clk),			// global clock input 
	.reset      (~reset_n),			// global reset input 

	.pbit       (cr_pbit),			// enable parity bit
	.ptype		(cr_ptype),			// type parity bit, 0 - even, 1 - odd
	.sbit       (cr_sbit),			// count stop bit, 2'b00 - 1 stop bit, 2'b01 - 2 stop bit, 2'b10 - 3 stop bit, 2'b11 - 3 stop bit;

	.ce_16      (ce_16),			// baud rate multiplyed by 16 - generated by baud module 
	.ser_in     (uart_rx),			// serial data input 
	
    .rx_data    (rx_data_o),		// data byte received 
	.new_rx_data(rx_valid_o),	// signs that a new byte was received 
	.pbit_error (rx_pbit_error)
);




endmodule